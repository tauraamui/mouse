module native

#include <linux/uinput.h>

struct C.uinput_setup {}

