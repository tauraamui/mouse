module main

import lib.display

fn main() {
	println(display.get_pixel_width_height())
}
